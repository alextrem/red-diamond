---------------------------------------
-- Company:
-- Engineer:        Alexander Geißler
--
-- Create Date:     23:40:00 02/26/2015
-- Design Name:
-- Project Name:    red-diamond
-- Target Device:   EP4CE22C8N
-- Tool Versions:   14.0
-- Description:     Audio interface of
-- ADV7612
--
-- Dependencies:
--
-- Revision:
-- Revision 0.1 - File created
--------------------------------------

